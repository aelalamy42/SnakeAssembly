library ieee; use ieee.std_logic_1164.all; use ieee.numeric_std.all; ENTiTy ID_S_B88a4C5_7E3415Ff_e is PORt( id_s_b88665f_7e7082e6_E : IN stD_LoGIC; iD_S_59777b_7ffcE7Ec_E : iN StD_lOgIc; id_s_16sgdbnv7_2c8dh7vjdo_E : In std_loGiC; id_s_c89sdnc7u_sda09scah_E : in std_lOgIc; iD_S_1F2653EB_6eC5B6Be_E : iN sTD_LoGic_vECtoR( 9 DOwnto 0); Id_S_25Bc52e8_112eF888_e : IN stD_logiC_VECtoR(31 DOwnTO 0); ID_S_191530B5_24e2b0bf_e : oUt StD_Logic_vEctoR(31 DOWNTo 0)); END ID_S_B88a4C5_7e3415fF_E; ArchitEcTUre ID_s_10643F3B_2fc543eB_E Of iD_s_B88A4C5_7e3415fF_E Is tyPe Id_S_77AfF7E5_27e78A14_E is aRRAY (0 To 1023) oF STd_lOgiC_vECtoR(31 dOWNTO 0); sIgNAL Id_S_B889004_7e48Ff67_e : id_S_77aFf7E5_27e78a14_e; signaL ID_S_cC3eE48_281C1fb9_E : Std_lOGic_vEctoR(9 DOwNTO 0); SignaL Id_S_6f8bcBE_62E8365d_e : sTd_lOgic; bEgIN ProCeSS(ID_s_B88665f_7e7082E6_E) bEgin if (Rising_edge(id_s_b88665F_7e7082e6_E) ) THen ID_S_6F8bcbE_62e8365D_E <= Id_s_59777B_7fFce7ec_E anD id_s_16sgdbnv7_2c8dh7vjdo_E; iD_s_cC3eE48_281c1fB9_E <= Id_s_1F2653eb_6eC5b6bE_E; eND IF; End PROCesS; Process(id_S_b889004_7e48FF67_E, ID_S_6F8bcBE_62E8365d_E, iD_s_CC3ee48_281C1FB9_E) BeGIn ID_S_191530B5_24E2B0Bf_E <= (others => 'Z'); IF (iD_s_6F8bCBE_62e8365D_E = '1') tHEN ID_S_191530B5_24e2B0BF_E <= ID_s_B889004_7e48fF67_E(To_IntegeR(UNsIgNeD(id_S_cC3ee48_281C1fb9_E))); END If; ENd prOceSS; PROcess(Id_S_B88665f_7E7082E6_e) bEgIn if (RiSiNG_edGe(ID_s_B88665F_7e7082E6_E) ) then if (id_s_59777b_7ffcE7EC_E = '1' AND id_s_c89sdnc7u_sda09scah_E = '1') then Id_s_B889004_7e48FF67_E( tO_INtEger(UNSigneD(id_s_1F2653eB_6eC5b6BE_E))) <= id_s_25Bc52E8_112EF888_E; eND IF; ENd If; enD PRoCeSs; EnD Id_s_10643F3B_2fC543eB_e;