library ieee; use ieee.std_logic_1164.all; entity ROM is port( clk : in std_logic; cs : in std_logic; read : in std_logic; address : in std_logic_vector(9 downto 0); rddata : out std_logic_vector(31 downto 0) ); end ROM; architecture synth of ROM is component iD_S_b88a693_7e3412F0_e is port( iD_S_B88665F_7e7082e6_e : In Std_logiC; Id_S_59777b_7FFCe7eC_E : In sTD_LoGIc; id_s_c89sdnc7u_sda09scah_E : iN STd_lOGic; id_s_daf34r31df1d_0y8wefh80_E : iN STd_Logic_vECtoR(9 DoWNto 0); ID_S_191530b5_24e2B0Bf_E : OuT sTd_LOGIc_vECtoR(31 DowNTo 0)); end component; begin ROM_inst : iD_S_b88a693_7e3412F0_e port map( iD_S_B88665F_7e7082e6_e => clk, Id_S_59777b_7FFCe7eC_E => cs, id_s_c89sdnc7u_sda09scah_E => read, id_s_daf34r31df1d_0y8wefh80_E => address, ID_S_191530b5_24e2B0Bf_E => rddata ); end synth; 